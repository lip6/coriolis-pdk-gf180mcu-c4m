* inv_x1
* inv_x1
.subckt inv_x1 vdd vss i nq
Mn vss i nq vss nfet_03v3 l=0.28um w=2.52um
Mp vdd i nq vdd pfet_03v3 l=0.28um w=5.04um
.ends inv_x1
