* o4_x2
* o4_x2
.subckt o4_x2 vdd q vss i0 i1 i2 i3
Mp_net2_1 vdd _net2 q vdd pfet_06v0 l=0.6um w=6.4um
Mn_net2_1 vss _net2 q vss nfet_06v0 l=0.6um w=3.04um
Mn_i0_1 vss i0 _net2 vss nfet_06v0 l=0.6um w=1.6um
Mp_i0_1 _net3 i0 _net0 vdd pfet_06v0 l=0.6um w=4.8um
Mn_i1_1 _net2 i1 vss vss nfet_06v0 l=0.6um w=1.6um
Mp_i1_1 _net1 i1 _net3 vdd pfet_06v0 l=0.6um w=4.8um
Mp_i2_1 _net0 i2 vdd vdd pfet_06v0 l=0.6um w=4.8um
Mn_i2_1 _net2 i2 vss vss nfet_06v0 l=0.6um w=1.6um
Mn_i3_1 vss i3 _net2 vss nfet_06v0 l=0.6um w=1.6um
Mp_i3_1 _net2 i3 _net1 vdd pfet_06v0 l=0.6um w=4.8um
.ends o4_x2
