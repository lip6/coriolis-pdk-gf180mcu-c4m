/*                                                                      */
/*  Avertec Release v3.4p5 (64 bits on Linux 5.4.109+)                  */
/*  [AVT_only] host: runner-xxurkrix-project-41071638-concurrent-0      */
/*  [AVT_only] arch: x86_64                                             */
/*  [AVT_only] path: /opt/tasyag-3.4p5/bin/avt_shell                    */
/*  argv:                                                               */
/*                                                                      */
/*  User: root                                                          */
/*  Generation date Mon May 22 11:35:14 2023                            */
/*                                                                      */
/*  Verilog data flow description generated from `sff1_x4`              */
/*                                                                      */


`timescale 1 ps/1 ps

module sff1_x4 (ck, i, q);

  input  ck;
  input  i;
  output q;

  reg sff_m;
  wire u;
  wire ck_delayed;

  assign ck'delayed = 1'bx;
  assign u = ~(i);

always @ (posedge ck)
begin
  sff_m <= ~(u);
end

  assign q = sff_m;

endmodule
