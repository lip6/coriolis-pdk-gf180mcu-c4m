* buf_x2
* buf_x2
.subckt buf_x2 vdd vss i q
Mn1 ni i vss vss nfet_06v0 l=0.6um w=1.6um
Mn2_0 vss ni q vss nfet_06v0 l=0.6um w=2.88um
Mn2_1 q ni vss vss nfet_06v0 l=0.6um w=2.88um
Mp1 ni i vdd vdd pfet_06v0 l=0.6um w=3.2um
Mp2_0 vdd ni q vdd pfet_06v0 l=0.6um w=5.76um
Mp2_1 q ni vdd vdd pfet_06v0 l=0.6um w=5.76um
.ends buf_x2
