* nand4_x0
.subckt nand4_x0 vdd vss nq i0 i1 i2 i3
Mn0 vss i0 int0 vss nfet_03v3 l=0.28um w=3.5um
Mp0 vdd i0 nq vdd pfet_03v3 l=0.28um w=3.5um
Mn1 int0 i1 int1 vss nfet_03v3 l=0.28um w=3.5um
Mp1 nq i1 vdd vdd pfet_03v3 l=0.28um w=3.5um
Mn2 int1 i2 int2 vss nfet_03v3 l=0.28um w=3.5um
Mp2 vdd i2 nq vdd pfet_03v3 l=0.28um w=3.5um
Mn3 int2 i3 nq vss nfet_03v3 l=0.28um w=3.5um
Mp3 nq i3 vdd vdd pfet_03v3 l=0.28um w=3.5um
.ends nand4_x0
