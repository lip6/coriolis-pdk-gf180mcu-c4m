* nxr2_x1
.subckt nxr2_x1 nq vdd vss i0 i1
Mp_net0_1 nq _net0 _net1 vdd pfet_03v3 l=0.28um w=5.6um
Mn_net0_1 nq _net0 _net2 vss nfet_03v3 l=0.28um w=2.66um
Mn_net3_1 _net4 _net3 nq vss nfet_03v3 l=0.28um w=2.66um
Mp_net3_1 _net1 _net3 vdd vdd pfet_03v3 l=0.28um w=5.6um
Mp_i0_1 _net0 i0 vdd vdd pfet_03v3 l=0.28um w=2.8um
Mn_i0_2 vss i0 _net4 vss nfet_03v3 l=0.28um w=2.66um
Mp_i0_2 vdd i0 _net1 vdd pfet_03v3 l=0.28um w=5.6um
Mn_i0_1 _net0 i0 vss vss nfet_03v3 l=0.28um w=1.4um
Mp_i1_1 _net1 i1 nq vdd pfet_03v3 l=0.28um w=5.6um
Mn_i1_1 _net2 i1 vss vss nfet_03v3 l=0.28um w=2.66um
Mp_i1_2 vdd i1 _net3 vdd pfet_03v3 l=0.28um w=2.8um
Mn_i1_2 vss i1 _net3 vss nfet_03v3 l=0.28um w=1.4um
.ends nxr2_x1
