* nxr2_x1
.subckt nxr2_x1 nq vdd vss i0 i1
Mp_net0_1 nq _net0 _net1 vdd pfet_06v0 l=0.6um w=6.4um
Mn_net0_1 nq _net0 _net2 vss nfet_06v0 l=0.6um w=3.04um
Mn_net3_1 _net4 _net3 nq vss nfet_06v0 l=0.6um w=3.04um
Mp_net3_1 _net1 _net3 vdd vdd pfet_06v0 l=0.6um w=6.4um
Mp_i0_1 _net0 i0 vdd vdd pfet_06v0 l=0.6um w=3.2um
Mn_i0_2 vss i0 _net4 vss nfet_06v0 l=0.6um w=3.04um
Mp_i0_2 vdd i0 _net1 vdd pfet_06v0 l=0.6um w=6.4um
Mn_i0_1 _net0 i0 vss vss nfet_06v0 l=0.6um w=1.6um
Mp_i1_1 _net1 i1 nq vdd pfet_06v0 l=0.6um w=6.4um
Mn_i1_1 _net2 i1 vss vss nfet_06v0 l=0.6um w=3.04um
Mp_i1_2 vdd i1 _net3 vdd pfet_06v0 l=0.6um w=3.2um
Mn_i1_2 vss i1 _net3 vss nfet_06v0 l=0.6um w=1.6um
.ends nxr2_x1
