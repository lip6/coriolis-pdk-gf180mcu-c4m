* one_x1
* one_x1
.subckt one_x1 vdd vss one
Mn vss one zero vss nfet_06v0 l=0.6um w=5.66um
Mp one zero vdd vdd pfet_06v0 l=0.6um w=6.3um
.ends one_x1
