* zeroone_x1
* zeroone_x1
.subckt zeroone_x1 vdd vss zero one
Mn vss one zero vss nfet_03v3 l=0.28um w=4.7um
Mp one zero vdd vdd pfet_03v3 l=0.28um w=5.26um
.ends zeroone_x1
