* zero_x1
* zero_x1
.subckt zero_x1 vdd vss zero
Mn vss one zero vss nfet_06v0 l=0.6um w=5.66um
Mp one zero vdd vdd pfet_06v0 l=0.6um w=6.3um
.ends zero_x1
