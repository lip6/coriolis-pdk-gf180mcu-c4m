* oa22_x2
.subckt oa22_x2 vdd q vss i0 i1 i2
Mp_net0_1 vdd _net0 q vdd pfet_03v3 l=0.28um w=5.6um
Mn_net0_1 vss _net0 q vss nfet_03v3 l=0.28um w=2.66um
Mn_i0_1 vss i0 _net2 vss nfet_03v3 l=0.28um w=2.66um
Mp_i0_1 _net1 i0 _net0 vdd pfet_03v3 l=0.28um w=2.8um
Mn_i1_1 _net2 i1 _net0 vss nfet_03v3 l=0.28um w=2.66um
Mp_i1_1 _net0 i1 _net1 vdd pfet_03v3 l=0.28um w=2.8um
Mp_i2_1 _net1 i2 vdd vdd pfet_03v3 l=0.28um w=2.8um
Mn_i2_1 _net0 i2 vss vss nfet_03v3 l=0.28um w=2.66um
.ends oa22_x2
