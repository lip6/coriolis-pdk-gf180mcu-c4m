* nand3_x0
.subckt nand3_x0 vdd vss nq i0 i1 i2
Mn0 vss i0 int0 vss nfet_06v0 l=0.6um w=4.0um
Mp0 vdd i0 nq vdd pfet_06v0 l=0.6um w=4.0um
Mn1 int0 i1 int1 vss nfet_06v0 l=0.6um w=4.0um
Mp1 nq i1 vdd vdd pfet_06v0 l=0.6um w=4.0um
Mn2 int1 i2 nq vss nfet_06v0 l=0.6um w=4.0um
Mp2 vdd i2 nq vdd pfet_06v0 l=0.6um w=4.0um
.ends nand3_x0
