* nor2_x0
* nor2_x0
.subckt nor2_x0 vdd vss nq i0 i1
Mn0 vss i0 nq vss nfet_03v3 l=0.28um w=1.4um
Mp0 vdd i0 int0 vdd pfet_03v3 l=0.28um w=4.2um
Mn1 nq i1 vss vss nfet_03v3 l=0.28um w=1.4um
Mp1 int0 i1 nq vdd pfet_03v3 l=0.28um w=4.2um
.ends nor2_x0
