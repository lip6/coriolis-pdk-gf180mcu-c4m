* a4_x2
* a4_x2
.subckt a4_x2 vdd q vss i0 i1 i2 i3
Mp_net1_1 vdd _net1 q vdd pfet_06v0 l=0.6um w=6.4um
Mn_net1_1 vss _net1 q vss nfet_06v0 l=0.6um w=3.04um
Mp_i0_1 vdd i0 _net1 vdd pfet_06v0 l=0.6um w=3.2um
Mn_i0_1 _net1 i0 _net3 vss nfet_06v0 l=0.6um w=3.2um
Mp_i1_1 _net1 i1 vdd vdd pfet_06v0 l=0.6um w=3.2um
Mn_i1_1 _net3 i1 _net0 vss nfet_06v0 l=0.6um w=3.2um
Mp_i2_1 vdd i2 _net1 vdd pfet_06v0 l=0.6um w=3.2um
Mn_i2_1 _net0 i2 _net2 vss nfet_06v0 l=0.6um w=3.2um
Mp_i3_1 _net1 i3 vdd vdd pfet_06v0 l=0.6um w=3.2um
Mn_i3_1 _net2 i3 vss vss nfet_06v0 l=0.6um w=3.2um
.ends a4_x2
