* a4_x2
* a4_x2
.subckt a4_x2 vdd q vss i0 i1 i2 i3
Mp_net1_1 vdd _net1 q vdd pfet_03v3 l=0.28um w=5.6um
Mn_net1_1 vss _net1 q vss nfet_03v3 l=0.28um w=2.66um
Mp_i0_1 vdd i0 _net1 vdd pfet_03v3 l=0.28um w=2.8um
Mn_i0_1 _net1 i0 _net3 vss nfet_03v3 l=0.28um w=2.8um
Mp_i1_1 _net1 i1 vdd vdd pfet_03v3 l=0.28um w=2.8um
Mn_i1_1 _net3 i1 _net0 vss nfet_03v3 l=0.28um w=2.8um
Mp_i2_1 vdd i2 _net1 vdd pfet_03v3 l=0.28um w=2.8um
Mn_i2_1 _net0 i2 _net2 vss nfet_03v3 l=0.28um w=2.8um
Mp_i3_1 _net1 i3 vdd vdd pfet_03v3 l=0.28um w=2.8um
Mn_i3_1 _net2 i3 vss vss nfet_03v3 l=0.28um w=2.8um
.ends a4_x2
