* a2_x2
* a2_x2
.subckt a2_x2 vss q vdd i0 i1
Mn_net0_1 vss _net0 q vss nfet_06v0 l=0.6um w=3.04um
Mp_net0_1 vdd _net0 q vdd pfet_06v0 l=0.6um w=6.4um
Mn_i0_1 _net0 i0 _net1 vss nfet_06v0 l=0.6um w=3.04um
Mp_i0_1 vdd i0 _net0 vdd pfet_06v0 l=0.6um w=3.2um
Mp_i1_1 _net0 i1 vdd vdd pfet_06v0 l=0.6um w=3.2um
Mn_i1_1 _net1 i1 vss vss nfet_06v0 l=0.6um w=3.04um
.ends a2_x2
