* nand2_x0
.subckt nand2_x0 vdd vss nq i0 i1
Mn0 vss i0 int0 vss nfet_03v3 l=0.28um w=2.8um
Mp0 vdd i0 nq vdd pfet_03v3 l=0.28um w=2.8um
Mn1 int0 i1 nq vss nfet_03v3 l=0.28um w=2.8um
Mp1 nq i1 vdd vdd pfet_03v3 l=0.28um w=2.8um
.ends nand2_x0
